module main

import vlibsql
import os

fn main() {
	env_path := '${@VMODROOT}/.env'
	load_env(env_path, false)
	libsql_url := os.getenv('LIBSQL_URL') or { panic('LIBSQL_URL not set in ${env_path}') }
	libsql_auth_token := os.getenv('LIBSQL_AUTH_TOKEN') or { panic('LIBSQL_AUTH_TOKEN not set in ${env_path}') }
	vlibsql.setup(vlibsql.Libsql_config_t{}) or { panic(err) }

	db := vlibsql.connect(
		url:        libsql_url
		path:       'local.db'
		auth_token: libsql_auth_token
	) or { panic(err) }

	defer {
		unsafe {
			db.free()
		}
	}

	setup_sql := "
	DROP TABLE IF EXISTS users;
	CREATE TABLE users (id INTEGER PRIMARY KEY AUTOINCREMENT, name TEXT);
	INSERT INTO users (name) VALUES ('Iku Turso');
	"
	db.batch(setup_sql) or { panic(err) }
	forenames := ['John', 'Jane', 'Jack', 'Jill']
	surnames := ['Smith', 'Doe', 'Black', 'White']

	mut stmt := db.prepare('INSERT INTO users (name) VALUES (?)') or { panic(err) }
	defer {
		unsafe {
			stmt.free()
		}
	}
	for forename in forenames {
		for surname in surnames {
			fullname := forename + ' ' + surname
			stmt.reset()
			stmt.bind_value(vlibsql.text(fullname)) or { panic(err) }
			stmt.execute() or { panic(err) }
		}
	}

	query_stmt := db.prepare('SELECT * FROM users') or { panic(err) }
	defer {
		unsafe {
			query_stmt.free()
		}
	}

	rows := query_stmt.query() or { panic(err) }
	for row in rows {
		id_ptr := row.value(0) or { panic(err) }
		name_ptr := row.value(1) or { panic(err) }
		unsafe {
			id := id_ptr.value.integer
			name := name_ptr.value.text.ptr
			println('id: ${id}')
			println('name: ${cstring_to_vstring(name)}')
		}
	}
}

fn load_env(path string, overwrite bool) {
	str := os.read_lines(path) or { panic(err) }
	for line in str {
		// Skip empty lines and comments
		env := line.split('=')
		key := env[0]
		value := env[1]
		os.setenv(key, value, overwrite)
	}
}
